`define DEFAULTSHARES 5
