`define DEFAULTSHARES 2
