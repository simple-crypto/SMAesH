localparam KSIZE_128 = 0;
localparam KSIZE_192 = 1;
localparam KSIZE_256 = 2;
