`define DEFAULTSHARES 3
