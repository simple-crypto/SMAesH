`define DEFAULTSHARES 4
